LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Trial_12 IS
GENERIC(SQUARE_HEIGHT : INTEGER := 50;
        SQUARE_WIDTH  : INTEGER := 50;
		  IM_WIDTH      : INTEGER := 55;  -- WIDTH  OF IMAGE1 IN MEMORY
        IM_HEIGHT     : INTEGER := 55;  -- HEIGHT OF IMAGE1 IN MEMORY
		  IM_WIDTH_1    : INTEGER := 200; -- WIDTH  OF IMAGE2 IN MEMORY
        IM_HEIGHT_1   : INTEGER := 133; -- HEIGHT OF IMAGE2 IN MEMORY
        DATASIZE      : INTEGER := 11;  -- MSB OF EACH ROW IN MEMORY
        ADDRESSSIZE   : INTEGER := 11;  -- MSB OF ADDRESSES
		  DATASIZE_2    : INTEGER := 11;  -- MSB OF EACH ROW IN MEMORY
        ADDRESSSIZE_2 : INTEGER := 14   -- MSB OF ADDRESSES
		  );

PORT(CLK50MHZ  : IN  STD_LOGIC;
	  KEY       : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
	  SW        : IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
	  LEDR      : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
     R         : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
     G         : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
     B         : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	  HEX0      : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	  HEX1      : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	  HEX2      : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
  	  HEX3      : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
     HSYNC     : OUT STD_LOGIC;
     VSYNC     : OUT STD_LOGIC);
END ENTITY Trial_12;

ARCHITECTURE DISPLAY OF Trial_12 IS
	-- PARAMETERS FOR A 1024X768 DISPLAY
	CONSTANT HFP768P  : INTEGER   := 24;
	CONSTANT HSP768P  : INTEGER   := 136;
	CONSTANT HBP768P  : INTEGER   := 160;
	CONSTANT HVA768P  : INTEGER   := 1024;
	CONSTANT HCN768P  : INTEGER   := 832;
	CONSTANT VFP768P  : INTEGER   := 3;
	CONSTANT VSP768P  : INTEGER   := 6;
	CONSTANT VBP768P  : INTEGER   := 29;
	CONSTANT VVA768P  : INTEGER   := 768;
	CONSTANT VCN768P  : INTEGER   := 422;
	CONSTANT VEN768P  : INTEGER   := 700;
	CONSTANT VTO768P  : INTEGER   := 100;
	CONSTANT VT1768P  : INTEGER   := 250;
	-- SIGNALS THAT WILL HOLD THE FRONT PORT ETC THAT WE WILL ACUTALLY USE
	SIGNAL   HFP      : INTEGER; -- HORIZONTAL FRONT PORCH
	SIGNAL   HSP      : INTEGER; -- HORIZONTAL SYNC PULSE
	SIGNAL   HBP      : INTEGER; -- HORIZONTAL BACK PORCH
	SIGNAL   HVA      : INTEGER; -- HORIZONTAL VISIBLE AREA
	SIGNAL   VFP      : INTEGER; -- VERTICAL FRONT PORCH
	SIGNAL   VSP      : INTEGER; -- VERTICAL SYNC PULSE
	SIGNAL   VBP      : INTEGER; -- VERTICAL BACK PORCH
	SIGNAL   VVA      : INTEGER; -- VERTICAL VISIBLE AREA
	SIGNAL   HCENTRE  : INTEGER;
	SIGNAL   VCENTRE  : INTEGER;
	SIGNAL   VEND     : INTEGER;
	SIGNAL   VTOP     : INTEGER;
	SIGNAL   VTOP1    : INTEGER;
	SIGNAL   START_P  : INTEGER;
	-- SIGNAL TO HOLD THE CLOCK WE WILL USE FOR THE DISPLAY
	SIGNAL  SYNC2_CLK : STD_LOGIC := '0';
	SIGNAL  SYNC_2CLK : STD_LOGIC := '0';
	SIGNAL  SW_CLK    : STD_LOGIC := '0';
	SIGNAL  P_CLK     : STD_LOGIC := '0';
	-- SIGNALS FOR EACH OF THE CLOCKS AVAILABLE TO US
	SIGNAL  CLK3_sec   : STD_LOGIC := '0';
	SIGNAL  CLK65      : STD_LOGIC := '0';
	SIGNAL  CLK_switch : STD_LOGIC := '0';
	SIGNAL  CLK_Play : STD_LOGIC := '0';
	-- SIGNALS TO HOLD THE PRESENT HORIZONTAL AND VERTICAL POSITIONS.
	SIGNAL HPOSITION  : INTEGER   := 0;
	SIGNAL VPOSITION  : INTEGER   := 0;
	-- SIGNALS TO HOLD THE PRESENT MEMORY ADDRESS TO BE READ AND THE DATA READ
	SIGNAL DATA_ADDRESS : STD_LOGIC_VECTOR(ADDRESSSIZE DOWNTO 0)   := (OTHERS=>'0');
	SIGNAL RAW_DATA     : STD_LOGIC_VECTOR(DATASIZE DOWNTO 0)      := (OTHERS=>'0');
	SIGNAL RAW_DATA_1   : STD_LOGIC_VECTOR(DATASIZE DOWNTO 0)      := (OTHERS=>'0');
	-- SIGNALS TO HOLD THE PRESENT MEMORY ADDRESS TO BE READ AND THE DATA READ
	SIGNAL DATA_ADDRESS_2 : STD_LOGIC_VECTOR(ADDRESSSIZE_2 DOWNTO 0)   := (OTHERS=>'0');
	SIGNAL RAW_DATA_2     : STD_LOGIC_VECTOR(DATASIZE_2 DOWNTO 0)      := (OTHERS=>'0');
	SIGNAL RAW_DATA_3     : STD_LOGIC_VECTOR(DATASIZE_2 DOWNTO 0)      := (OTHERS=>'0');
	-- SIGNALS TO HOLD IMAGE DIMESIONS
	SIGNAL IMAGE1_HEIGHT  : INTEGER   := 0;
	SIGNAL IMAGE1_WIDTH   : INTEGER   := 0;
	-- SIGNALS TO HOLD IMAGE DIMESIONS
	SIGNAL IMAGE2_HEIGHT  : INTEGER   := 0;
	SIGNAL IMAGE2_WIDTH   : INTEGER   := 0;

	
	SIGNAL Dir, Ri                   : STD_LOGIC;
	SIGNAL SHOOT                              : STD_LOGIC := '1';
	SIGNAL KILL                               : STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL K1, K2, K3, K4, K5, K6             : STD_LOGIC := '0';
	SIGNAL SWITCH                             : STD_LOGIC := '1';
	SIGNAL U                                  : STD_LOGIC := '0';
	SIGNAL W                                  : STD_LOGIC := '0';
	SIGNAL V                                  : STD_LOGIC := '0';
	SIGNAL F                                  : STD_LOGIC_VECTOR(1 DOWNTO 0):=    "00";
	SIGNAL P                                  : STD_LOGIC_VECTOR(5 DOWNTO 0):="000000"; --VARIABLE TO COMPARE TO KILL
	
	
BEGIN
	SYNC_2CLK <= CLK3_sec;
	SYNC2_CLK <= CLK65;
	SW_CLK    <= CLK_switch;
	P_CLK     <= CLK_play;
	HFP       <= HFP768P;
	HSP       <= HSP768P;
	HBP       <= HBP768P;
	HVA       <= HVA768P;
	VFP       <= VFP768P;
	VSP       <= VSP768P;
	VBP       <= VBP768P;
	VVA       <= VVA768P;
	HCENTRE   <= HCN768P;
	VCENTRE   <= VCN768P;
	VEND      <= VEN768P;
	VTOP      <= VTO768P;
	VTOP1     <= VT1768P;
	IMAGE1_HEIGHT <=   IM_HEIGHT;
	IMAGE1_WIDTH  <=    IM_WIDTH;
	IMAGE2_HEIGHT <= IM_HEIGHT_1;
	IMAGE2_WIDTH  <=  IM_WIDTH_1;
	Ri  <= KEY(0);
	Dir <= SW(0);
	
	LEDR(9) <= U;
	LEDR(8) <= W;
	
	DISP_CLK:   WORK.sec_3_clk    PORT MAP(clk_1  => CLK50MHZ,
										         T0     => CLK3_sec);
	DISP_CLK_1: WORK.CLK_SYNQ     PORT MAP(INCLK0 => CLK50MHZ,
												   C0     => CLK65);
	DISP_CLK_2: WORK.switch_clk   PORT MAP(clk_2 => CLK50MHZ,
												   T1     => CLK_switch);
	DISP_CLK_3: WORK.Pl_CLK       PORT MAP(clk_3 => CLK50MHZ,
												   T2     => CLK_play);
	IMRED:		WORK.IMREAD       PORT MAP(ADDRESS => DATA_ADDRESS,
													CLOCK    => SYNC2_CLK,
													Q        => RAW_DATA);
	IMRED_1:    WORK.IMREAD_1     PORT MAP(ADDRESS => DATA_ADDRESS,
												   CLOCK    => SYNC2_CLK,
													Q        => RAW_DATA_1);
	IMRED_2:    WORK.IMREAD_2     PORT MAP(ADDRESS => DATA_ADDRESS_2,
												   CLOCK    => SYNC2_CLK,
													Q        => RAW_DATA_2);
	IMRED_3:    WORK.IMREAD_3     PORT MAP(ADDRESS => DATA_ADDRESS_2,
												   CLOCK    => SYNC2_CLK,
													Q        => RAW_DATA_3);
	
	PROCESS(SYNC2_CLK, SYNC_2CLK, SW_CLK, P_CLK, Ri, SWITCH, U, V, W, Dir, K6, K5, K4, K3, K2, K1, P, KILL, F)
	
	VARIABLE START_P  : INTEGER := 800;
	VARIABLE START_E1 : INTEGER := 700;
	VARIABLE START_E2 : INTEGER := 800;
	VARIABLE START_E3 : INTEGER := 900;
	VARIABLE START_E4 : INTEGER := 700;
	VARIABLE START_E5 : INTEGER := 800;
	VARIABLE START_E6 : INTEGER := 900;
	VARIABLE END_HSTART          : INTEGER := 500;
	VARIABLE END_HSTOP           : INTEGER := END_HSTART + IMAGE2_WIDTH;
	VARIABLE END_VSTART          : INTEGER := 500;
	VARIABLE END_VSTOP           : INTEGER := END_VSTART + IMAGE2_HEIGHT;
	VARIABLE IMAGE1_HSTART       : INTEGER := START_E1;
	VARIABLE IMAGE1_HSTOP        : INTEGER := IMAGE1_HSTART + IMAGE1_WIDTH;
	VARIABLE IMAGE1_VSTART       : INTEGER := VTOP;
	VARIABLE IMAGE1_VSTOP        : INTEGER := IMAGE1_VSTART + IMAGE1_HEIGHT;
	VARIABLE IMAGE2_HSTART       : INTEGER := START_E2;
	VARIABLE IMAGE2_HSTOP        : INTEGER := IMAGE2_HSTART + IMAGE1_WIDTH;
	VARIABLE IMAGE2_VSTART       : INTEGER := VTOP;
	VARIABLE IMAGE2_VSTOP        : INTEGER := IMAGE2_VSTART + IMAGE1_HEIGHT;
	VARIABLE IMAGE3_HSTART       : INTEGER := START_E3;
	VARIABLE IMAGE3_HSTOP        : INTEGER := IMAGE3_HSTART + IMAGE1_WIDTH;
	VARIABLE IMAGE3_VSTART       : INTEGER := VTOP;
	VARIABLE IMAGE3_VSTOP        : INTEGER := IMAGE3_VSTART + IMAGE1_HEIGHT;
	VARIABLE IMAGE4_HSTART       : INTEGER := START_E4;
	VARIABLE IMAGE4_HSTOP        : INTEGER := IMAGE4_HSTART + IMAGE1_WIDTH;
	VARIABLE IMAGE4_VSTART       : INTEGER := VTOP1;
	VARIABLE IMAGE4_VSTOP        : INTEGER := IMAGE4_VSTART + IMAGE1_HEIGHT;
	VARIABLE IMAGE5_HSTART       : INTEGER := START_E5;
	VARIABLE IMAGE5_HSTOP        : INTEGER := IMAGE5_HSTART + IMAGE1_WIDTH;
	VARIABLE IMAGE5_VSTART       : INTEGER := VTOP1;
	VARIABLE IMAGE5_VSTOP        : INTEGER := IMAGE5_VSTART + IMAGE1_HEIGHT;
	VARIABLE IMAGE6_HSTART       : INTEGER := START_E6;
	VARIABLE IMAGE6_HSTOP        : INTEGER := IMAGE6_HSTART + IMAGE1_WIDTH;
	VARIABLE IMAGE6_VSTART       : INTEGER := VTOP1;
	VARIABLE IMAGE6_VSTOP        : INTEGER := IMAGE6_VSTART + IMAGE1_HEIGHT;
	
	VARIABLE IMAGE1_PIXEL_COL, IMAGE1_PIXEL_ROW, IMAGE1_PIXEL_NUMBER    : INTEGER := 0;
	VARIABLE IMAGE2_PIXEL_COL, IMAGE2_PIXEL_ROW, IMAGE2_PIXEL_NUMBER    : INTEGER := 0;
	VARIABLE IMAGE3_PIXEL_COL, IMAGE3_PIXEL_ROW, IMAGE3_PIXEL_NUMBER    : INTEGER := 0;
	VARIABLE IMAGE4_PIXEL_COL, IMAGE4_PIXEL_ROW, IMAGE4_PIXEL_NUMBER    : INTEGER := 0;
	VARIABLE IMAGE5_PIXEL_COL, IMAGE5_PIXEL_ROW, IMAGE5_PIXEL_NUMBER    : INTEGER := 0;
	VARIABLE IMAGE6_PIXEL_COL, IMAGE6_PIXEL_ROW, IMAGE6_PIXEL_NUMBER    : INTEGER := 0;
	VARIABLE END_PIXEL_COL   , END_PIXEL_ROW   , END_PIXEL_NUMBER       : INTEGER := 0;
	VARIABLE B_POS              : INTEGER := 650;
	VARIABLE START_B            : INTEGER :=   0;
	VARIABLE MEM_ADDRESS        : UNSIGNED(ADDRESSSIZE   DOWNTO 0) := (OTHERS=>'0');
	VARIABLE MEM_ADDRESS_2      : UNSIGNED(ADDRESSSIZE_2 DOWNTO 0) := (OTHERS=>'0');
	
	VARIABLE K_COUNT : INTEGER := 0; -- VARIABLE TO HOLD KILL COUNT
	VARIABLE N       : INTEGER := 0; -- VARIABLE TO COMPARE TO SHOTT
	
	BEGIN

		KILL  <= K6 & K5 & K4 & K3 & K2 & K1;
				
		IF Ri <= '0' THEN
			SHOOT <= '0';
		ELSIF Ri <= '1' THEN
			SHOOT <= '1';
		END IF;
		
		IF RISING_EDGE(Ri) THEN
			N := N + 1;
		END IF;
		
		IF N = 10 AND K_COUNT < 6 THEN
			F <= "10";
		ELSIF N > 10 AND K_COUNT < 6 THEN
			F <= "10";
		ELSIF K_COUNT = 6 THEN
			F <= "01";
		ELSE
			F <= "00";
		END IF;
		
		IF RISING_EDGE(SYNC_2CLK) THEN
			
			LEDR(0)          <=       SHOOT;
			
			IF SHOOT <= '0' THEN
				B_POS := B_POS - 20;
			ELSIF SHOOT <= '1' THEN
				B_POS := 650;
			END IF;
			
			IF (START_E1 < 400) THEN
				U <= '0';
			ELSIF START_E3 > 1200 THEN
				U <= '1';
			END IF;
			
			IF (START_E4 < 400) THEN
				W <= '1';
			ELSIF START_E6 > 1200 THEN
				W <= '0';
			END IF;
			
			IF P = KILL THEN
				K_COUNT := K_COUNT;
			ELSIF P /= KILL THEN
				K_COUNT := K_COUNT + 1;
				P <= KILL;
			END IF;
			
			IF K_COUNT = 0 THEN
				HEX2 <= STD_LOGIC_VECTOR'("01000000");
				HEX3 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF K_COUNT = 1 THEN
				HEX2 <= STD_LOGIC_VECTOR'("01111001");
				HEX3 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF K_COUNT = 2 THEN
				HEX2 <= STD_LOGIC_VECTOR'("00100100");
				HEX3 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF K_COUNT = 3 THEN
				HEX2 <= STD_LOGIC_VECTOR'("00110000");
				HEX3 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF K_COUNT = 4 THEN
				HEX2 <= STD_LOGIC_VECTOR'("00011001");
				HEX3 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF K_COUNT = 5 THEN
				HEX2 <= STD_LOGIC_VECTOR'("00010010");
				HEX3 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF K_COUNT = 6 THEN
				HEX2 <= STD_LOGIC_VECTOR'("00000010");
				HEX3 <= STD_LOGIC_VECTOR'("11000000");
			ELSE
				HEX2 <= STD_LOGIC_VECTOR'("11111111");
				HEX3 <= STD_LOGIC_VECTOR'("11111111");
			END IF;
			
			IF N = 0 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF N = 1 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF N = 2 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF N = 3 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF N = 4 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF N = 5 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF N = 6 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF N = 7 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF N = 8 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF N = 9 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF N = 10 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSE
				HEX0 <= STD_LOGIC_VECTOR'("11111111");
				HEX1 <= STD_LOGIC_VECTOR'("11111111");
			END IF;
			
			IF U <= '0' THEN
				START_E1 := START_E1 + 40;
				START_E2 := START_E2 + 40;
				START_E3 := START_E3 + 40;
			ELSIF U <= '1' THEN
				START_E1 := START_E1 - 40;
				START_E2 := START_E2 - 40;
				START_E3 := START_E3 - 40;
			END IF;	
				
			IF W <= '0' THEN	
				START_E4 := START_E4 - 40;
				START_E5 := START_E5 - 40;
				START_E6 := START_E6 - 40;
			ELSIF W <= '1' THEN
				START_E4 := START_E4 + 40;
				START_E5 := START_E5 + 40;
				START_E6 := START_E6 + 40;
			END IF;
				
			IF (B_POS > 100) AND (B_POS < 155) THEN
				IF (START_B > IMAGE1_HSTART) AND (START_B < IMAGE1_HSTOP) THEN
					K1 <= '1';
				ELSIF (START_B > IMAGE2_HSTART) AND (START_B < IMAGE2_HSTOP) THEN
					K2 <= '1';
				ELSIF (START_B > IMAGE3_HSTART) AND (START_B < IMAGE3_HSTOP) THEN
					K3 <= '1';
				END IF;
			ELSIF (B_POS > 250) AND (B_POS < 305) THEN
				IF (START_B > IMAGE4_HSTART) AND (START_B < IMAGE4_HSTOP) THEN
					K4 <= '1';
				ELSIF (START_B > IMAGE5_HSTART) AND (START_B < IMAGE5_HSTOP) THEN
					K5 <= '1';
				ELSIF (START_B > IMAGE6_HSTART) AND (START_B < IMAGE6_HSTOP) THEN
					K6 <= '1';
				END IF;
			END IF;
		END IF;
		
		IF RISING_EDGE(P_CLK) THEN
		
			IF (START_P < 450) THEN
				V <= '0';
			ELSIF START_P > 1200 THEN
				V <= '1';
			ELSIF Dir = '0' THEN
				V <= '1';
			ELSIF Dir = '1' THEN
				V <= '0';
			END IF;
			
			IF V <= '0' THEN
				START_P := START_P + 40;
			ELSIF V <= '1' THEN
				START_P := START_P - 40;
			END IF;
		END IF;
			
		IF RISING_EDGE(SW_CLK) THEN
			SWITCH <= NOT(SWITCH);
		END IF;
			
		IF RISING_EDGE(SYNC2_CLK) THEN
			-- ALWAYS INCREMENT THE HORIZONTAL POSITION COUNTER WITH EACH ACTIVE CLOCK PULSE
			HPOSITION <= HPOSITION + 1;
			
			-- WHEN HORIZONTAL POSITION COUNTER GETS TO THE LAST PIXEL IN A ROW, GO BACK
			-- TO ZERO AND INCREMENT THE VERTICAL COUNTER (I.E. GO TO START OF NEXT LINE)
			IF HPOSITION >= (HFP+HSP+HBP+HVA) THEN
				HPOSITION <= 0;
				-- WHEN VERTICAL POSITION COUNTER GETS TO THE END OF ROWS, GO BACK TO THE
				-- START OF THE FIRST ROW
				IF VPOSITION >= (VFP+VSP+VBP+VVA) THEN
					VPOSITION <= 0;
				ELSE
					VPOSITION <= VPOSITION + 1;
				END IF;
			END IF;
			
			
			-- GENERATE HORIZONTAL SYNCH PULSE WHENEVER THE HPOSITION IS BETWEEN THE FRONT
			-- PORCH AND THE BACK PORCH
			IF (HPOSITION >= HFP) AND (HPOSITION < (HFP+HSP)) THEN
				HSYNC <= '0';
			ELSE
				HSYNC <= '1';
			END IF;
			
			-- GENERATE VERTICAL SYNCH PULSE WHENEVER THE VPOSITION IS BETWEEN THE FRONT
			-- PORCH AND THE BACK PORCH
			IF (VPOSITION >= VFP) AND (VPOSITION < (VFP+VSP)) THEN
				VSYNC <= '0';
			ELSE
				VSYNC <= '1';
			END IF;
			
			
			-- NOW TO PUT THINGS UP ON THE DISPLAY
			-- WHERE DO WE WANT TO PUT THINGS?
			-- LET'S PUT THE IMAGE IN OUR MEMORY IN THE CENTRE OF THE SCREEN STARTING
			-- FROM THE 100TH ROW. WE FIRST DETERMINE THE BOUNDS IN WHICH THE IMAGE WILL BE
			-- DISPLAYED AND THEN TELL IT WHAT MEMORY ADDRESS TO READ FROM IN ORDER TO 
			-- DISPLAY THE CONTENTS OF THE MEMORY ONTO THE DISPLAY.
			-- THE CENTRAL PIXEL OF THE VISIBLE AREA IS 
			
			IF F = "00" THEN
			
				IF SHOOT <= '0' THEN
									
					IF START_B = 0 THEN
						START_B := START_P;
					ELSE
						START_B := START_B;
					END IF;
						
					IF (VPOSITION > (B_POS) AND VPOSITION <= (B_POS + 20)) AND (HPOSITION >= (START_B - 3) AND HPOSITION <= (START_B + 3)) THEN
						R <= X"F";
						G <= X"0";
						B <= X"0";
					ELSIF (VPOSITION > VEND AND VPOSITION <= (VEND + (SQUARE_HEIGHT/2))) AND (HPOSITION >= (START_P - (SQUARE_WIDTH/4)) AND HPOSITION <= (START_P + (SQUARE_WIDTH/4))) THEN
						R <= X"A";
						G <= X"1";
						B <= X"7";
					ELSIF (VPOSITION > (VEND + (SQUARE_HEIGHT/2)) AND VPOSITION <= (VEND + SQUARE_HEIGHT)) AND (HPOSITION >= (START_P - (SQUARE_WIDTH)) AND HPOSITION <= (START_P + (SQUARE_WIDTH))) THEN
						R <= X"F";
						G <= X"1";
						B <= X"1";
					ELSIF (HPOSITION >= IMAGE1_HSTART AND HPOSITION <= IMAGE1_HSTOP) AND (VPOSITION >= IMAGE1_VSTART AND VPOSITION <= IMAGE1_VSTOP) THEN
						IF K1 <= '0' THEN
							IMAGE1_PIXEL_COL := HPOSITION - IMAGE1_HSTART;
							IMAGE1_PIXEL_ROW := VPOSITION - IMAGE1_VSTART;
							IMAGE1_PIXEL_NUMBER := IMAGE1_PIXEL_COL + IMAGE1_PIXEL_ROW*IMAGE1_WIDTH;
							MEM_ADDRESS  := TO_UNSIGNED(IMAGE1_PIXEL_NUMBER, MEM_ADDRESS'LENGTH);
							DATA_ADDRESS <= STD_LOGIC_VECTOR(MEM_ADDRESS);
							IF SWITCH <= '0' THEN
								R <= RAW_DATA(11 DOWNTO 8);
								G <= RAW_DATA(7 DOWNTO 4);
								B <= RAW_DATA(3 DOWNTO 0);
							ELSE
								R <= RAW_DATA_1(11 DOWNTO 8);
								G <= RAW_DATA_1(7 DOWNTO 4);
								B <= RAW_DATA_1(3 DOWNTO 0);
							END IF;
						ELSE
							R <= X"0";
							G <= X"0";
							B <= X"0";
						END IF;
					ELSIF (HPOSITION >= IMAGE2_HSTART AND HPOSITION <= IMAGE2_HSTOP) AND (VPOSITION >= IMAGE2_VSTART AND VPOSITION <= IMAGE2_VSTOP) THEN
						IF K2 <= '0' THEN	
							IMAGE2_PIXEL_COL := HPOSITION - IMAGE2_HSTART;
							IMAGE2_PIXEL_ROW := VPOSITION - IMAGE2_VSTART;
							IMAGE2_PIXEL_NUMBER := IMAGE2_PIXEL_COL + IMAGE2_PIXEL_ROW*IMAGE1_WIDTH;
							MEM_ADDRESS  := TO_UNSIGNED(IMAGE2_PIXEL_NUMBER, MEM_ADDRESS'LENGTH);
							DATA_ADDRESS <= STD_LOGIC_VECTOR(MEM_ADDRESS);
							IF SWITCH <= '0' THEN
								R <= RAW_DATA(11 DOWNTO 8);
								G <= RAW_DATA(7 DOWNTO 4);
								B <= RAW_DATA(3 DOWNTO 0);
							ELSE
								R <= RAW_DATA_1(11 DOWNTO 8);
								G <= RAW_DATA_1(7 DOWNTO 4);
								B <= RAW_DATA_1(3 DOWNTO 0);
							END IF;
						ELSE
							R <= X"0";
							G <= X"0";
							B <= X"0";
						END IF;
					ELSIF (HPOSITION >= IMAGE3_HSTART AND HPOSITION <= IMAGE3_HSTOP) AND (VPOSITION >= IMAGE3_VSTART AND VPOSITION <= IMAGE3_VSTOP) THEN
						IF K3 <= '0' THEN	
							IMAGE3_PIXEL_COL := HPOSITION - IMAGE3_HSTART;
							IMAGE3_PIXEL_ROW := VPOSITION - IMAGE3_VSTART;
							IMAGE3_PIXEL_NUMBER := IMAGE3_PIXEL_COL + IMAGE3_PIXEL_ROW*IMAGE1_WIDTH;
							MEM_ADDRESS  := TO_UNSIGNED(IMAGE3_PIXEL_NUMBER, MEM_ADDRESS'LENGTH);
							DATA_ADDRESS <= STD_LOGIC_VECTOR(MEM_ADDRESS);
							IF SWITCH <= '0' THEN
								R <= RAW_DATA(11 DOWNTO 8);
								G <= RAW_DATA(7 DOWNTO 4);
								B <= RAW_DATA(3 DOWNTO 0);
							ELSE
								R <= RAW_DATA_1(11 DOWNTO 8);
								G <= RAW_DATA_1(7 DOWNTO 4);
								B <= RAW_DATA_1(3 DOWNTO 0);
							END IF;
						ELSE
							R <= X"0";
							G <= X"0";
							B <= X"0";
						END IF;
					ELSIF (HPOSITION >= IMAGE4_HSTART AND HPOSITION <= IMAGE4_HSTOP) AND (VPOSITION >= IMAGE4_VSTART AND VPOSITION <= IMAGE4_VSTOP) THEN
						IF K4 <= '0' THEN	
							IMAGE4_PIXEL_COL := HPOSITION - IMAGE4_HSTART;
							IMAGE4_PIXEL_ROW := VPOSITION - IMAGE4_VSTART;
							IMAGE4_PIXEL_NUMBER := IMAGE4_PIXEL_COL + IMAGE4_PIXEL_ROW*IMAGE1_WIDTH;
							MEM_ADDRESS  := TO_UNSIGNED(IMAGE4_PIXEL_NUMBER, MEM_ADDRESS'LENGTH);
							DATA_ADDRESS <= STD_LOGIC_VECTOR(MEM_ADDRESS);
							IF SWITCH <= '0' THEN
								R <= RAW_DATA(11 DOWNTO 8);
								G <= RAW_DATA(7 DOWNTO 4);
								B <= RAW_DATA(3 DOWNTO 0);
							ELSE
								R <= RAW_DATA_1(11 DOWNTO 8);
								G <= RAW_DATA_1(7 DOWNTO 4);
								B <= RAW_DATA_1(3 DOWNTO 0);
							END IF;
						ELSE
							R <= X"0";
							G <= X"0";
							B <= X"0";
						END IF;
					ELSIF (HPOSITION >= IMAGE5_HSTART AND HPOSITION <= IMAGE5_HSTOP) AND (VPOSITION >= IMAGE5_VSTART AND VPOSITION <= IMAGE5_VSTOP) THEN
						IF K5 <= '0' THEN	
							IMAGE5_PIXEL_COL := HPOSITION - IMAGE5_HSTART;
							IMAGE5_PIXEL_ROW := VPOSITION - IMAGE5_VSTART;
							IMAGE5_PIXEL_NUMBER := IMAGE5_PIXEL_COL + IMAGE5_PIXEL_ROW*IMAGE1_WIDTH;
							MEM_ADDRESS  := TO_UNSIGNED(IMAGE5_PIXEL_NUMBER, MEM_ADDRESS'LENGTH);
							DATA_ADDRESS <= STD_LOGIC_VECTOR(MEM_ADDRESS);
							IF SWITCH <= '0' THEN
								R <= RAW_DATA(11 DOWNTO 8);
								G <= RAW_DATA(7 DOWNTO 4);
								B <= RAW_DATA(3 DOWNTO 0);
							ELSE
								R <= RAW_DATA_1(11 DOWNTO 8);
								G <= RAW_DATA_1(7 DOWNTO 4);
								B <= RAW_DATA_1(3 DOWNTO 0);
							END IF;
						ELSE
							R <= X"0";
							G <= X"0";
							B <= X"0";
						END IF;
					ELSIF (HPOSITION >= IMAGE6_HSTART AND HPOSITION <= IMAGE6_HSTOP) AND (VPOSITION >= IMAGE6_VSTART AND VPOSITION <= IMAGE6_VSTOP) THEN
						IF K6 <= '0' THEN	
							IMAGE6_PIXEL_COL := HPOSITION - IMAGE6_HSTART;
							IMAGE6_PIXEL_ROW := VPOSITION - IMAGE6_VSTART;
							IMAGE6_PIXEL_NUMBER := IMAGE6_PIXEL_COL + IMAGE6_PIXEL_ROW*IMAGE1_WIDTH;
							MEM_ADDRESS  := TO_UNSIGNED(IMAGE6_PIXEL_NUMBER, MEM_ADDRESS'LENGTH);
							DATA_ADDRESS <= STD_LOGIC_VECTOR(MEM_ADDRESS);
							IF SWITCH <= '0' THEN
								R <= RAW_DATA(11 DOWNTO 8);
								G <= RAW_DATA(7 DOWNTO 4);
								B <= RAW_DATA(3 DOWNTO 0);
							ELSE
								R <= RAW_DATA_1(11 DOWNTO 8);
								G <= RAW_DATA_1(7 DOWNTO 4);
								B <= RAW_DATA_1(3 DOWNTO 0);
							END IF;
						ELSE
							R <= X"0";
							G <= X"0";
							B <= X"0";
						END IF;
					ELSE
						R <= X"0";
						G <= X"0";
						B <= X"0";
					END IF;
				ELSE
					
					START_B := 0;
					
					IF (VPOSITION > VEND AND VPOSITION <= (VEND + (SQUARE_HEIGHT/2))) AND (HPOSITION >= (START_P - (SQUARE_WIDTH/4)) AND HPOSITION <= (START_P + (SQUARE_WIDTH/4))) THEN
						R <= X"A";
						G <= X"1";
						B <= X"7";
					ELSIF (VPOSITION > (VEND + (SQUARE_HEIGHT/2)) AND VPOSITION <= (VEND + SQUARE_HEIGHT)) AND (HPOSITION >= (START_P - (SQUARE_WIDTH)) AND HPOSITION <= (START_P + (SQUARE_WIDTH))) THEN
						R <= X"7";
						G <= X"1";
						B <= X"A";
					ELSIF (HPOSITION >= IMAGE1_HSTART AND HPOSITION <= IMAGE1_HSTOP) AND (VPOSITION >= IMAGE1_VSTART AND VPOSITION <= IMAGE1_VSTOP) THEN
						IF K1 <= '0' THEN
							IMAGE1_PIXEL_COL := HPOSITION - IMAGE1_HSTART;
							IMAGE1_PIXEL_ROW := VPOSITION - IMAGE1_VSTART;
							IMAGE1_PIXEL_NUMBER := IMAGE1_PIXEL_COL + IMAGE1_PIXEL_ROW*IMAGE1_WIDTH;
							MEM_ADDRESS  := TO_UNSIGNED(IMAGE1_PIXEL_NUMBER, MEM_ADDRESS'LENGTH);
							DATA_ADDRESS <= STD_LOGIC_VECTOR(MEM_ADDRESS);
							IF SWITCH <= '0' THEN
								R <= RAW_DATA(11 DOWNTO 8);
								G <= RAW_DATA(7 DOWNTO 4);
								B <= RAW_DATA(3 DOWNTO 0);
							ELSE
								R <= RAW_DATA_1(11 DOWNTO 8);
								G <= RAW_DATA_1(7 DOWNTO 4);
								B <= RAW_DATA_1(3 DOWNTO 0);
							END IF;
						ELSE
							R <= X"0";
							G <= X"0";
							B <= X"0";
						END IF;
					ELSIF (HPOSITION >= IMAGE2_HSTART AND HPOSITION <= IMAGE2_HSTOP) AND (VPOSITION >= IMAGE2_VSTART AND VPOSITION <= IMAGE2_VSTOP) THEN
						IF K2 <= '0' THEN	
							IMAGE2_PIXEL_COL := HPOSITION - IMAGE2_HSTART;
							IMAGE2_PIXEL_ROW := VPOSITION - IMAGE2_VSTART;
							IMAGE2_PIXEL_NUMBER := IMAGE2_PIXEL_COL + IMAGE2_PIXEL_ROW*IMAGE1_WIDTH;
							MEM_ADDRESS  := TO_UNSIGNED(IMAGE2_PIXEL_NUMBER, MEM_ADDRESS'LENGTH);
							DATA_ADDRESS <= STD_LOGIC_VECTOR(MEM_ADDRESS);
							IF SWITCH <= '0' THEN
								R <= RAW_DATA(11 DOWNTO 8);
								G <= RAW_DATA(7 DOWNTO 4);
								B <= RAW_DATA(3 DOWNTO 0);
							ELSE
								R <= RAW_DATA_1(11 DOWNTO 8);
								G <= RAW_DATA_1(7 DOWNTO 4);
								B <= RAW_DATA_1(3 DOWNTO 0);
							END IF;
						ELSE
							R <= X"0";
							G <= X"0";
							B <= X"0";
						END IF;
					ELSIF (HPOSITION >= IMAGE3_HSTART AND HPOSITION <= IMAGE3_HSTOP) AND (VPOSITION >= IMAGE3_VSTART AND VPOSITION <= IMAGE3_VSTOP) THEN
						IF K3 <= '0' THEN	
							IMAGE3_PIXEL_COL := HPOSITION - IMAGE3_HSTART;
							IMAGE3_PIXEL_ROW := VPOSITION - IMAGE3_VSTART;
							IMAGE3_PIXEL_NUMBER := IMAGE3_PIXEL_COL + IMAGE3_PIXEL_ROW*IMAGE1_WIDTH;
							MEM_ADDRESS  := TO_UNSIGNED(IMAGE3_PIXEL_NUMBER, MEM_ADDRESS'LENGTH);
							DATA_ADDRESS <= STD_LOGIC_VECTOR(MEM_ADDRESS);
							IF SWITCH <= '0' THEN
								R <= RAW_DATA(11 DOWNTO 8);
								G <= RAW_DATA(7 DOWNTO 4);
								B <= RAW_DATA(3 DOWNTO 0);
							ELSE
								R <= RAW_DATA_1(11 DOWNTO 8);
								G <= RAW_DATA_1(7 DOWNTO 4);
								B <= RAW_DATA_1(3 DOWNTO 0);
							END IF;
						ELSE
							R <= X"0";
							G <= X"0";
							B <= X"0";
						END IF;
					ELSIF (HPOSITION >= IMAGE4_HSTART AND HPOSITION <= IMAGE4_HSTOP) AND (VPOSITION >= IMAGE4_VSTART AND VPOSITION <= IMAGE4_VSTOP) THEN
						IF K4 <= '0' THEN	
							IMAGE4_PIXEL_COL := HPOSITION - IMAGE4_HSTART;
							IMAGE4_PIXEL_ROW := VPOSITION - IMAGE4_VSTART;
							IMAGE4_PIXEL_NUMBER := IMAGE4_PIXEL_COL + IMAGE4_PIXEL_ROW*IMAGE1_WIDTH;
							MEM_ADDRESS  := TO_UNSIGNED(IMAGE4_PIXEL_NUMBER, MEM_ADDRESS'LENGTH);
							DATA_ADDRESS <= STD_LOGIC_VECTOR(MEM_ADDRESS);
							IF SWITCH <= '0' THEN
								R <= RAW_DATA(11 DOWNTO 8);
								G <= RAW_DATA(7 DOWNTO 4);
								B <= RAW_DATA(3 DOWNTO 0);
							ELSE
								R <= RAW_DATA_1(11 DOWNTO 8);
								G <= RAW_DATA_1(7 DOWNTO 4);
								B <= RAW_DATA_1(3 DOWNTO 0);
							END IF;
						ELSE
							R <= X"0";
							G <= X"0";
							B <= X"0";
						END IF;
					ELSIF (HPOSITION >= IMAGE5_HSTART AND HPOSITION <= IMAGE5_HSTOP) AND (VPOSITION >= IMAGE5_VSTART AND VPOSITION <= IMAGE5_VSTOP) THEN
						IF K5 <= '0' THEN	
							IMAGE5_PIXEL_COL := HPOSITION - IMAGE5_HSTART;
							IMAGE5_PIXEL_ROW := VPOSITION - IMAGE5_VSTART;
							IMAGE5_PIXEL_NUMBER := IMAGE5_PIXEL_COL + IMAGE5_PIXEL_ROW*IMAGE1_WIDTH;
							MEM_ADDRESS  := TO_UNSIGNED(IMAGE5_PIXEL_NUMBER, MEM_ADDRESS'LENGTH);
							DATA_ADDRESS <= STD_LOGIC_VECTOR(MEM_ADDRESS);
							IF SWITCH <= '0' THEN
								R <= RAW_DATA(11 DOWNTO 8);
								G <= RAW_DATA(7 DOWNTO 4);
								B <= RAW_DATA(3 DOWNTO 0);
							ELSE
								R <= RAW_DATA_1(11 DOWNTO 8);
								G <= RAW_DATA_1(7 DOWNTO 4);
								B <= RAW_DATA_1(3 DOWNTO 0);
							END IF;
						ELSE
							R <= X"0";
							G <= X"0";
							B <= X"0";
						END IF;
					ELSIF (HPOSITION >= IMAGE6_HSTART AND HPOSITION <= IMAGE6_HSTOP) AND (VPOSITION >= IMAGE6_VSTART AND VPOSITION <= IMAGE6_VSTOP) THEN
						IF K6 <= '0' THEN	
							IMAGE6_PIXEL_COL := HPOSITION - IMAGE6_HSTART;
							IMAGE6_PIXEL_ROW := VPOSITION - IMAGE6_VSTART;
							IMAGE6_PIXEL_NUMBER := IMAGE6_PIXEL_COL + IMAGE6_PIXEL_ROW*IMAGE1_WIDTH;
							MEM_ADDRESS  := TO_UNSIGNED(IMAGE6_PIXEL_NUMBER, MEM_ADDRESS'LENGTH);
							DATA_ADDRESS <= STD_LOGIC_VECTOR(MEM_ADDRESS);
							IF SWITCH <= '0' THEN
								R <= RAW_DATA(11 DOWNTO 8);
								G <= RAW_DATA(7 DOWNTO 4);
								B <= RAW_DATA(3 DOWNTO 0);
							ELSE
								R <= RAW_DATA_1(11 DOWNTO 8);
								G <= RAW_DATA_1(7 DOWNTO 4);
								B <= RAW_DATA_1(3 DOWNTO 0);
							END IF;
						ELSE
							R <= X"0";
							G <= X"0";
							B <= X"0";
						END IF;
					ELSE
						R <= X"0";
						G <= X"0";
						B <= X"0";
					END IF;
				END IF;
			ELSIF F = "01" THEN
				IF (HPOSITION >= (HCENTRE - (IMAGE2_WIDTH/2)) AND HPOSITION <= (HCENTRE + (IMAGE2_WIDTH/2))) AND (VPOSITION >= (VCENTRE - (IMAGE2_HEIGHT/2)) AND VPOSITION <= (VCENTRE + (IMAGE2_HEIGHT/2))) THEN
					END_PIXEL_COL := HPOSITION - END_HSTART;
					END_PIXEL_ROW := VPOSITION - END_VSTART;
					END_PIXEL_NUMBER := END_PIXEL_COL + END_PIXEL_ROW*IMAGE2_WIDTH;
					MEM_ADDRESS_2  := TO_UNSIGNED(END_PIXEL_NUMBER, MEM_ADDRESS_2'LENGTH);
					DATA_ADDRESS_2 <= STD_LOGIC_VECTOR(MEM_ADDRESS_2);
						R <= RAW_DATA_2(11 DOWNTO 8);
						G <= RAW_DATA_2(7 DOWNTO 4);
						B <= RAW_DATA_2(3 DOWNTO 0);
				ELSE
					R <= X"0";
					G <= X"0";
					B <= X"0";
				END IF;
			ELSIF F = "10" THEN
				IF (HPOSITION >= (HCENTRE - (IMAGE2_WIDTH/2)) AND HPOSITION <= (HCENTRE + (IMAGE2_WIDTH/2))) AND (VPOSITION >= (VCENTRE - (IMAGE2_HEIGHT/2)) AND VPOSITION <= (VCENTRE + (IMAGE2_HEIGHT/2))) THEN
					END_PIXEL_COL := HPOSITION - END_HSTART;
					END_PIXEL_ROW := VPOSITION - END_VSTART;
					END_PIXEL_NUMBER := END_PIXEL_COL + END_PIXEL_ROW*IMAGE2_WIDTH;
					MEM_ADDRESS_2  := TO_UNSIGNED(END_PIXEL_NUMBER, MEM_ADDRESS_2'LENGTH);
					DATA_ADDRESS_2 <= STD_LOGIC_VECTOR(MEM_ADDRESS_2);
						R <= RAW_DATA_3(11 DOWNTO 8);
						G <= RAW_DATA_3(7 DOWNTO 4);
						B <= RAW_DATA_3(3 DOWNTO 0);
				ELSE
					R <= X"0";
					G <= X"0";
					B <= X"0";
				END IF;
			END IF;
		END IF;
	END PROCESS;

END ARCHITECTURE DISPLAY;